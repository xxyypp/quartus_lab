count8_inst : count8 PORT MAP (
		clock	 => clock_sig,
		q	 => q_sig
	);
