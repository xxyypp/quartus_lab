flip_inst : flip PORT MAP (
		clock	 => clock_sig,
		q	 => q_sig
	);
